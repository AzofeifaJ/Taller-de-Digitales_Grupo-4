module ImgROM (
    input   wire            i_clk,
    input   wire            i_res_n,
    input   wire    [12:0]  i_addr,
    output  reg     [ 7:0]  o_data
    );
    always @(posedge i_clk or negedge i_res_n) begin
        if (~i_res_n) begin
            o_data <= 8'd0;
        end else begin
            o_data <= imageROM( i_addr );
        end
    end
    
    function [7:0] imageROM;
        input   [12:0]   addr;
        begin
            case (addr)
                0: imageROM = 8'd63;
                1: imageROM = 8'd63;
                2: imageROM = 8'd63;
                3: imageROM = 8'd63;
                4: imageROM = 8'd63;
                5: imageROM = 8'd63;
                6: imageROM = 8'd63;
                7: imageROM = 8'd63;
                8: imageROM = 8'd63;
                9: imageROM = 8'd63;
                10: imageROM = 8'd63;
                11: imageROM = 8'd63;
                12: imageROM = 8'd63;
                13: imageROM = 8'd63;
                14: imageROM = 8'd63;
                15: imageROM = 8'd25;
                16: imageROM = 8'd77;
                17: imageROM = 8'd63;
                18: imageROM = 8'd47;
                19: imageROM = 8'd88;
                20: imageROM = 8'd63;
                21: imageROM = 8'd38;
                22: imageROM = 8'd94;
                23: imageROM = 8'd63;
                24: imageROM = 8'd33;
                25: imageROM = 8'd98;
                26: imageROM = 8'd63;
                27: imageROM = 8'd29;
                28: imageROM = 8'd102;
                29: imageROM = 8'd63;
                30: imageROM = 8'd25;
                31: imageROM = 8'd106;
                32: imageROM = 8'd63;
                33: imageROM = 8'd21;
                34: imageROM = 8'd78;
                35: imageROM = 8'd146;
                36: imageROM = 8'd77;
                37: imageROM = 8'd63;
                38: imageROM = 8'd18;
                39: imageROM = 8'd76;
                40: imageROM = 8'd154;
                41: imageROM = 8'd74;
                42: imageROM = 8'd63;
                43: imageROM = 8'd16;
                44: imageROM = 8'd75;
                45: imageROM = 8'd158;
                46: imageROM = 8'd73;
                47: imageROM = 8'd63;
                48: imageROM = 8'd14;
                49: imageROM = 8'd73;
                50: imageROM = 8'd163;
                51: imageROM = 8'd72;
                52: imageROM = 8'd63;
                53: imageROM = 8'd12;
                54: imageROM = 8'd73;
                55: imageROM = 8'd165;
                56: imageROM = 8'd72;
                57: imageROM = 8'd63;
                58: imageROM = 8'd10;
                59: imageROM = 8'd72;
                60: imageROM = 8'd168;
                61: imageROM = 8'd72;
                62: imageROM = 8'd63;
                63: imageROM = 8'd8;
                64: imageROM = 8'd72;
                65: imageROM = 8'd171;
                66: imageROM = 8'd71;
                67: imageROM = 8'd63;
                68: imageROM = 8'd6;
                69: imageROM = 8'd71;
                70: imageROM = 8'd135;
                71: imageROM = 8'd69;
                72: imageROM = 8'd161;
                73: imageROM = 8'd71;
                74: imageROM = 8'd63;
                75: imageROM = 8'd5;
                76: imageROM = 8'd71;
                77: imageROM = 8'd135;
                78: imageROM = 8'd71;
                79: imageROM = 8'd159;
                80: imageROM = 8'd73;
                81: imageROM = 8'd63;
                82: imageROM = 8'd3;
                83: imageROM = 8'd71;
                84: imageROM = 8'd135;
                85: imageROM = 8'd73;
                86: imageROM = 8'd141;
                87: imageROM = 8'd72;
                88: imageROM = 8'd136;
                89: imageROM = 8'd74;
                90: imageROM = 8'd63;
                91: imageROM = 8'd2;
                92: imageROM = 8'd71;
                93: imageROM = 8'd136;
                94: imageROM = 8'd73;
                95: imageROM = 8'd139;
                96: imageROM = 8'd76;
                97: imageROM = 8'd134;
                98: imageROM = 8'd75;
                99: imageROM = 8'd63;
                100: imageROM = 8'd1;
                101: imageROM = 8'd70;
                102: imageROM = 8'd137;
                103: imageROM = 8'd74;
                104: imageROM = 8'd136;
                105: imageROM = 8'd79;
                106: imageROM = 8'd133;
                107: imageROM = 8'd75;
                108: imageROM = 8'd63;
                109: imageROM = 8'd70;
                110: imageROM = 8'd138;
                111: imageROM = 8'd74;
                112: imageROM = 8'd135;
                113: imageROM = 8'd81;
                114: imageROM = 8'd132;
                115: imageROM = 8'd76;
                116: imageROM = 8'd61;
                117: imageROM = 8'd71;
                118: imageROM = 8'd138;
                119: imageROM = 8'd74;
                120: imageROM = 8'd135;
                121: imageROM = 8'd82;
                122: imageROM = 8'd131;
                123: imageROM = 8'd76;
                124: imageROM = 8'd61;
                125: imageROM = 8'd70;
                126: imageROM = 8'd139;
                127: imageROM = 8'd74;
                128: imageROM = 8'd134;
                129: imageROM = 8'd84;
                130: imageROM = 8'd130;
                131: imageROM = 8'd77;
                132: imageROM = 8'd59;
                133: imageROM = 8'd70;
                134: imageROM = 8'd140;
                135: imageROM = 8'd74;
                136: imageROM = 8'd134;
                137: imageROM = 8'd70;
                138: imageROM = 8'd199;
                139: imageROM = 8'd71;
                140: imageROM = 8'd130;
                141: imageROM = 8'd77;
                142: imageROM = 8'd59;
                143: imageROM = 8'd70;
                144: imageROM = 8'd140;
                145: imageROM = 8'd74;
                146: imageROM = 8'd133;
                147: imageROM = 8'd71;
                148: imageROM = 8'd200;
                149: imageROM = 8'd71;
                150: imageROM = 8'd130;
                151: imageROM = 8'd76;
                152: imageROM = 8'd58;
                153: imageROM = 8'd70;
                154: imageROM = 8'd142;
                155: imageROM = 8'd73;
                156: imageROM = 8'd133;
                157: imageROM = 8'd70;
                158: imageROM = 8'd202;
                159: imageROM = 8'd70;
                160: imageROM = 8'd131;
                161: imageROM = 8'd69;
                162: imageROM = 8'd129;
                163: imageROM = 8'd70;
                164: imageROM = 8'd57;
                165: imageROM = 8'd70;
                166: imageROM = 8'd143;
                167: imageROM = 8'd71;
                168: imageROM = 8'd134;
                169: imageROM = 8'd70;
                170: imageROM = 8'd202;
                171: imageROM = 8'd70;
                172: imageROM = 8'd133;
                173: imageROM = 8'd66;
                174: imageROM = 8'd130;
                175: imageROM = 8'd70;
                176: imageROM = 8'd57;
                177: imageROM = 8'd70;
                178: imageROM = 8'd144;
                179: imageROM = 8'd69;
                180: imageROM = 8'd134;
                181: imageROM = 8'd70;
                182: imageROM = 8'd204;
                183: imageROM = 8'd70;
                184: imageROM = 8'd137;
                185: imageROM = 8'd70;
                186: imageROM = 8'd55;
                187: imageROM = 8'd70;
                188: imageROM = 8'd156;
                189: imageROM = 8'd70;
                190: imageROM = 8'd204;
                191: imageROM = 8'd70;
                192: imageROM = 8'd137;
                193: imageROM = 8'd70;
                194: imageROM = 8'd55;
                195: imageROM = 8'd70;
                196: imageROM = 8'd156;
                197: imageROM = 8'd70;
                198: imageROM = 8'd204;
                199: imageROM = 8'd70;
                200: imageROM = 8'd138;
                201: imageROM = 8'd70;
                202: imageROM = 8'd54;
                203: imageROM = 8'd69;
                204: imageROM = 8'd157;
                205: imageROM = 8'd70;
                206: imageROM = 8'd204;
                207: imageROM = 8'd70;
                208: imageROM = 8'd139;
                209: imageROM = 8'd69;
                210: imageROM = 8'd53;
                211: imageROM = 8'd70;
                212: imageROM = 8'd157;
                213: imageROM = 8'd70;
                214: imageROM = 8'd205;
                215: imageROM = 8'd69;
                216: imageROM = 8'd139;
                217: imageROM = 8'd70;
                218: imageROM = 8'd52;
                219: imageROM = 8'd70;
                220: imageROM = 8'd157;
                221: imageROM = 8'd70;
                222: imageROM = 8'd205;
                223: imageROM = 8'd70;
                224: imageROM = 8'd138;
                225: imageROM = 8'd70;
                226: imageROM = 8'd52;
                227: imageROM = 8'd70;
                228: imageROM = 8'd156;
                229: imageROM = 8'd71;
                230: imageROM = 8'd205;
                231: imageROM = 8'd70;
                232: imageROM = 8'd139;
                233: imageROM = 8'd69;
                234: imageROM = 8'd52;
                235: imageROM = 8'd69;
                236: imageROM = 8'd158;
                237: imageROM = 8'd70;
                238: imageROM = 8'd205;
                239: imageROM = 8'd70;
                240: imageROM = 8'd139;
                241: imageROM = 8'd70;
                242: imageROM = 8'd50;
                243: imageROM = 8'd70;
                244: imageROM = 8'd158;
                245: imageROM = 8'd70;
                246: imageROM = 8'd205;
                247: imageROM = 8'd70;
                248: imageROM = 8'd139;
                249: imageROM = 8'd70;
                250: imageROM = 8'd50;
                251: imageROM = 8'd70;
                252: imageROM = 8'd158;
                253: imageROM = 8'd70;
                254: imageROM = 8'd205;
                255: imageROM = 8'd70;
                256: imageROM = 8'd139;
                257: imageROM = 8'd70;
                258: imageROM = 8'd50;
                259: imageROM = 8'd70;
                260: imageROM = 8'd158;
                261: imageROM = 8'd70;
                262: imageROM = 8'd205;
                263: imageROM = 8'd70;
                264: imageROM = 8'd140;
                265: imageROM = 8'd69;
                266: imageROM = 8'd50;
                267: imageROM = 8'd69;
                268: imageROM = 8'd159;
                269: imageROM = 8'd70;
                270: imageROM = 8'd205;
                271: imageROM = 8'd70;
                272: imageROM = 8'd140;
                273: imageROM = 8'd70;
                274: imageROM = 8'd48;
                275: imageROM = 8'd70;
                276: imageROM = 8'd159;
                277: imageROM = 8'd70;
                278: imageROM = 8'd205;
                279: imageROM = 8'd70;
                280: imageROM = 8'd140;
                281: imageROM = 8'd70;
                282: imageROM = 8'd48;
                283: imageROM = 8'd70;
                284: imageROM = 8'd159;
                285: imageROM = 8'd70;
                286: imageROM = 8'd205;
                287: imageROM = 8'd70;
                288: imageROM = 8'd140;
                289: imageROM = 8'd70;
                290: imageROM = 8'd47;
                291: imageROM = 8'd70;
                292: imageROM = 8'd161;
                293: imageROM = 8'd70;
                294: imageROM = 8'd204;
                295: imageROM = 8'd70;
                296: imageROM = 8'd141;
                297: imageROM = 8'd69;
                298: imageROM = 8'd47;
                299: imageROM = 8'd70;
                300: imageROM = 8'd161;
                301: imageROM = 8'd70;
                302: imageROM = 8'd203;
                303: imageROM = 8'd70;
                304: imageROM = 8'd142;
                305: imageROM = 8'd69;
                306: imageROM = 8'd47;
                307: imageROM = 8'd69;
                308: imageROM = 8'd162;
                309: imageROM = 8'd70;
                310: imageROM = 8'd203;
                311: imageROM = 8'd70;
                312: imageROM = 8'd142;
                313: imageROM = 8'd69;
                314: imageROM = 8'd46;
                315: imageROM = 8'd70;
                316: imageROM = 8'd162;
                317: imageROM = 8'd70;
                318: imageROM = 8'd203;
                319: imageROM = 8'd70;
                320: imageROM = 8'd142;
                321: imageROM = 8'd69;
                322: imageROM = 8'd46;
                323: imageROM = 8'd70;
                324: imageROM = 8'd163;
                325: imageROM = 8'd69;
                326: imageROM = 8'd203;
                327: imageROM = 8'd70;
                328: imageROM = 8'd142;
                329: imageROM = 8'd69;
                330: imageROM = 8'd45;
                331: imageROM = 8'd70;
                332: imageROM = 8'd164;
                333: imageROM = 8'd70;
                334: imageROM = 8'd201;
                335: imageROM = 8'd70;
                336: imageROM = 8'd143;
                337: imageROM = 8'd69;
                338: imageROM = 8'd45;
                339: imageROM = 8'd70;
                340: imageROM = 8'd164;
                341: imageROM = 8'd70;
                342: imageROM = 8'd201;
                343: imageROM = 8'd70;
                344: imageROM = 8'd142;
                345: imageROM = 8'd70;
                346: imageROM = 8'd44;
                347: imageROM = 8'd71;
                348: imageROM = 8'd165;
                349: imageROM = 8'd70;
                350: imageROM = 8'd199;
                351: imageROM = 8'd71;
                352: imageROM = 8'd142;
                353: imageROM = 8'd70;
                354: imageROM = 8'd44;
                355: imageROM = 8'd70;
                356: imageROM = 8'd166;
                357: imageROM = 8'd70;
                358: imageROM = 8'd198;
                359: imageROM = 8'd71;
                360: imageROM = 8'd143;
                361: imageROM = 8'd70;
                362: imageROM = 8'd43;
                363: imageROM = 8'd71;
                364: imageROM = 8'd166;
                365: imageROM = 8'd71;
                366: imageROM = 8'd197;
                367: imageROM = 8'd71;
                368: imageROM = 8'd143;
                369: imageROM = 8'd70;
                370: imageROM = 8'd43;
                371: imageROM = 8'd71;
                372: imageROM = 8'd167;
                373: imageROM = 8'd71;
                374: imageROM = 8'd195;
                375: imageROM = 8'd71;
                376: imageROM = 8'd144;
                377: imageROM = 8'd69;
                378: imageROM = 8'd43;
                379: imageROM = 8'd72;
                380: imageROM = 8'd168;
                381: imageROM = 8'd70;
                382: imageROM = 8'd195;
                383: imageROM = 8'd70;
                384: imageROM = 8'd144;
                385: imageROM = 8'd70;
                386: imageROM = 8'd43;
                387: imageROM = 8'd72;
                388: imageROM = 8'd168;
                389: imageROM = 8'd71;
                390: imageROM = 8'd193;
                391: imageROM = 8'd71;
                392: imageROM = 8'd144;
                393: imageROM = 8'd70;
                394: imageROM = 8'd42;
                395: imageROM = 8'd73;
                396: imageROM = 8'd169;
                397: imageROM = 8'd77;
                398: imageROM = 8'd145;
                399: imageROM = 8'd70;
                400: imageROM = 8'd41;
                401: imageROM = 8'd74;
                402: imageROM = 8'd170;
                403: imageROM = 8'd76;
                404: imageROM = 8'd145;
                405: imageROM = 8'd69;
                406: imageROM = 8'd42;
                407: imageROM = 8'd75;
                408: imageROM = 8'd170;
                409: imageROM = 8'd74;
                410: imageROM = 8'd145;
                411: imageROM = 8'd70;
                412: imageROM = 8'd41;
                413: imageROM = 8'd76;
                414: imageROM = 8'd170;
                415: imageROM = 8'd73;
                416: imageROM = 8'd146;
                417: imageROM = 8'd70;
                418: imageROM = 8'd41;
                419: imageROM = 8'd76;
                420: imageROM = 8'd171;
                421: imageROM = 8'd72;
                422: imageROM = 8'd146;
                423: imageROM = 8'd69;
                424: imageROM = 8'd41;
                425: imageROM = 8'd70;
                426: imageROM = 8'd130;
                427: imageROM = 8'd70;
                428: imageROM = 8'd171;
                429: imageROM = 8'd70;
                430: imageROM = 8'd146;
                431: imageROM = 8'd70;
                432: imageROM = 8'd40;
                433: imageROM = 8'd71;
                434: imageROM = 8'd130;
                435: imageROM = 8'd70;
                436: imageROM = 8'd171;
                437: imageROM = 8'd70;
                438: imageROM = 8'd146;
                439: imageROM = 8'd70;
                440: imageROM = 8'd39;
                441: imageROM = 8'd71;
                442: imageROM = 8'd132;
                443: imageROM = 8'd70;
                444: imageROM = 8'd171;
                445: imageROM = 8'd68;
                446: imageROM = 8'd146;
                447: imageROM = 8'd70;
                448: imageROM = 8'd40;
                449: imageROM = 8'd70;
                450: imageROM = 8'd133;
                451: imageROM = 8'd70;
                452: imageROM = 8'd172;
                453: imageROM = 8'd67;
                454: imageROM = 8'd146;
                455: imageROM = 8'd70;
                456: imageROM = 8'd39;
                457: imageROM = 8'd71;
                458: imageROM = 8'd134;
                459: imageROM = 8'd70;
                460: imageROM = 8'd191;
                461: imageROM = 8'd129;
                462: imageROM = 8'd70;
                463: imageROM = 8'd38;
                464: imageROM = 8'd71;
                465: imageROM = 8'd135;
                466: imageROM = 8'd71;
                467: imageROM = 8'd190;
                468: imageROM = 8'd70;
                469: imageROM = 8'd38;
                470: imageROM = 8'd71;
                471: imageROM = 8'd137;
                472: imageROM = 8'd70;
                473: imageROM = 8'd190;
                474: imageROM = 8'd70;
                475: imageROM = 8'd37;
                476: imageROM = 8'd71;
                477: imageROM = 8'd139;
                478: imageROM = 8'd70;
                479: imageROM = 8'd189;
                480: imageROM = 8'd69;
                481: imageROM = 8'd37;
                482: imageROM = 8'd71;
                483: imageROM = 8'd140;
                484: imageROM = 8'd71;
                485: imageROM = 8'd187;
                486: imageROM = 8'd70;
                487: imageROM = 8'd36;
                488: imageROM = 8'd72;
                489: imageROM = 8'd141;
                490: imageROM = 8'd71;
                491: imageROM = 8'd186;
                492: imageROM = 8'd70;
                493: imageROM = 8'd35;
                494: imageROM = 8'd72;
                495: imageROM = 8'd143;
                496: imageROM = 8'd71;
                497: imageROM = 8'd185;
                498: imageROM = 8'd69;
                499: imageROM = 8'd35;
                500: imageROM = 8'd72;
                501: imageROM = 8'd145;
                502: imageROM = 8'd72;
                503: imageROM = 8'd182;
                504: imageROM = 8'd70;
                505: imageROM = 8'd35;
                506: imageROM = 8'd71;
                507: imageROM = 8'd147;
                508: imageROM = 8'd72;
                509: imageROM = 8'd181;
                510: imageROM = 8'd70;
                511: imageROM = 8'd34;
                512: imageROM = 8'd71;
                513: imageROM = 8'd149;
                514: imageROM = 8'd73;
                515: imageROM = 8'd179;
                516: imageROM = 8'd69;
                517: imageROM = 8'd34;
                518: imageROM = 8'd71;
                519: imageROM = 8'd151;
                520: imageROM = 8'd74;
                521: imageROM = 8'd176;
                522: imageROM = 8'd70;
                523: imageROM = 8'd33;
                524: imageROM = 8'd71;
                525: imageROM = 8'd153;
                526: imageROM = 8'd77;
                527: imageROM = 8'd172;
                528: imageROM = 8'd70;
                529: imageROM = 8'd32;
                530: imageROM = 8'd71;
                531: imageROM = 8'd156;
                532: imageROM = 8'd82;
                533: imageROM = 8'd165;
                534: imageROM = 8'd70;
                535: imageROM = 8'd32;
                536: imageROM = 8'd71;
                537: imageROM = 8'd157;
                538: imageROM = 8'd81;
                539: imageROM = 8'd165;
                540: imageROM = 8'd70;
                541: imageROM = 8'd31;
                542: imageROM = 8'd71;
                543: imageROM = 8'd160;
                544: imageROM = 8'd79;
                545: imageROM = 8'd165;
                546: imageROM = 8'd70;
                547: imageROM = 8'd30;
                548: imageROM = 8'd71;
                549: imageROM = 8'd164;
                550: imageROM = 8'd76;
                551: imageROM = 8'd165;
                552: imageROM = 8'd70;
                553: imageROM = 8'd29;
                554: imageROM = 8'd71;
                555: imageROM = 8'd167;
                556: imageROM = 8'd74;
                557: imageROM = 8'd165;
                558: imageROM = 8'd69;
                559: imageROM = 8'd29;
                560: imageROM = 8'd71;
                561: imageROM = 8'd174;
                562: imageROM = 8'd66;
                563: imageROM = 8'd167;
                564: imageROM = 8'd69;
                565: imageROM = 8'd28;
                566: imageROM = 8'd71;
                567: imageROM = 8'd191;
                568: imageROM = 8'd153;
                569: imageROM = 8'd70;
                570: imageROM = 8'd26;
                571: imageROM = 8'd71;
                572: imageROM = 8'd191;
                573: imageROM = 8'd154;
                574: imageROM = 8'd70;
                575: imageROM = 8'd25;
                576: imageROM = 8'd71;
                577: imageROM = 8'd191;
                578: imageROM = 8'd155;
                579: imageROM = 8'd70;
                580: imageROM = 8'd24;
                581: imageROM = 8'd71;
                582: imageROM = 8'd191;
                583: imageROM = 8'd156;
                584: imageROM = 8'd70;
                585: imageROM = 8'd23;
                586: imageROM = 8'd71;
                587: imageROM = 8'd191;
                588: imageROM = 8'd157;
                589: imageROM = 8'd70;
                590: imageROM = 8'd22;
                591: imageROM = 8'd71;
                592: imageROM = 8'd191;
                593: imageROM = 8'd158;
                594: imageROM = 8'd70;
                595: imageROM = 8'd21;
                596: imageROM = 8'd71;
                597: imageROM = 8'd191;
                598: imageROM = 8'd160;
                599: imageROM = 8'd69;
                600: imageROM = 8'd20;
                601: imageROM = 8'd71;
                602: imageROM = 8'd191;
                603: imageROM = 8'd161;
                604: imageROM = 8'd70;
                605: imageROM = 8'd18;
                606: imageROM = 8'd71;
                607: imageROM = 8'd191;
                608: imageROM = 8'd162;
                609: imageROM = 8'd70;
                610: imageROM = 8'd18;
                611: imageROM = 8'd70;
                612: imageROM = 8'd191;
                613: imageROM = 8'd163;
                614: imageROM = 8'd70;
                615: imageROM = 8'd17;
                616: imageROM = 8'd70;
                617: imageROM = 8'd191;
                618: imageROM = 8'd165;
                619: imageROM = 8'd69;
                620: imageROM = 8'd17;
                621: imageROM = 8'd70;
                622: imageROM = 8'd191;
                623: imageROM = 8'd165;
                624: imageROM = 8'd70;
                625: imageROM = 8'd16;
                626: imageROM = 8'd69;
                627: imageROM = 8'd191;
                628: imageROM = 8'd167;
                629: imageROM = 8'd69;
            endcase
        end
    endfunction
endmodule